interface hvac_intf(input logic clk,reset);

logic I1;
logic I2;
logic I3;
logic I4;
logic O1;
logic O2;
logic O3;
logic O4;

endinterface

