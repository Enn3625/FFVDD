`include "usr.v"
`include "transaction.sv"
`include "generator.sv"
`include "hvac_intf.sv"
`include "bfm.sv"
`include "environment.sv"
`include "hvac_test.sv"
`include "top.sv"




